erik@erik-VirtualBox.20531:1435260824